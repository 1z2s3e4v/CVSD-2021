/home/raid7_1/userd/d10013/CVSD/lab6/Lab6/library/lef/tsmc13fsg_8lm_cic.lef