

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO ipdc 
  PIN i_clk 
    ANTENNAPARTIALMETALAREA 0.101 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3535 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 55.534 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 194.509 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 32.776 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 114.856 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0556 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 31.8585 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 111.221 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.102596 LAYER VIA45 ;
  END i_clk
  PIN i_rst_n 
    ANTENNAPARTIALMETALAREA 56.828 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 199.178 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2106 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 270.64 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 948.098 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAMAXCUTCAR 0.34283 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 17.324 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 61.194 LAYER METAL3 ;
    ANTENNAGATEAREA 2.2789 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 278.242 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 974.95 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.850078 LAYER VIA34 ;
  END i_rst_n
  PIN i_op_valid 
    ANTENNAPARTIALMETALAREA 54.733 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 191.566 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 2.58 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.31 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.065 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 87.6708 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 317.837 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 3.33231 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 1.162 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 4.207 LAYER METAL5 ;
    ANTENNAGATEAREA 0.1638 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 94.7648 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 343.521 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 3.33231 LAYER VIA56 ;
  END i_op_valid
  PIN i_op_mode[3] 
    ANTENNAPARTIALMETALAREA 55.662 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 194.957 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 2.436 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.666 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0988 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 48.1412 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 172.893 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.09615 LAYER VIA45 ;
  END i_op_mode[3]
  PIN i_op_mode[2] 
    ANTENNAPARTIALMETALAREA 55.662 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 194.957 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 2.62 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.31 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0845 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 37.8982 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 136.724 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.28166 LAYER VIA45 ;
  END i_op_mode[2]
  PIN i_op_mode[1] 
    ANTENNAPARTIALMETALAREA 57.722 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 202.167 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.334 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.309 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1157 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 19.9801 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 70.8712 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.624028 LAYER VIA34 ;
  END i_op_mode[1]
  PIN i_op_mode[0] 
    ANTENNAPARTIALMETALAREA 59.396 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 207.886 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1157 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 519.157 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 1815.06 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.312014 LAYER VIA23 ;
  END i_op_mode[0]
  PIN o_op_ready 
    ANTENNADIFFAREA 0.7208 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 59.844 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 209.594 LAYER METAL2 ;
  END o_op_ready
  PIN i_in_valid 
    ANTENNAPARTIALMETALAREA 65.204 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 228.354 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3458 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 191.345 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 667.772 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.514245 LAYER VIA23 ;
  END i_in_valid
  PIN i_in_data[23] 
    ANTENNAPARTIALMETALAREA 21.092 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 73.822 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 20.758 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 72.793 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL5 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA56 ;
    ANTENNAPARTIALMETALAREA 30.48 LAYER METAL6 ;
    ANTENNAPARTIALMETALSIDEAREA 106.82 LAYER METAL6 ;
  END i_in_data[23]
  PIN i_in_data[22] 
    ANTENNAPARTIALMETALAREA 20.764 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 72.674 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 10.27 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 36.085 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL5 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA56 ;
    ANTENNAPARTIALMETALAREA 30.972 LAYER METAL6 ;
    ANTENNAPARTIALMETALSIDEAREA 108.542 LAYER METAL6 ;
  END i_in_data[22]
  PIN i_in_data[21] 
    ANTENNAPARTIALMETALAREA 18.786 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 65.751 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.334 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.309 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL5 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA56 ;
    ANTENNAPARTIALMETALAREA 32.612 LAYER METAL6 ;
    ANTENNAPARTIALMETALSIDEAREA 114.282 LAYER METAL6 ;
  END i_in_data[21]
  PIN i_in_data[20] 
    ANTENNAPARTIALMETALAREA 81.8706 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 285.947 LAYER METAL2 ;
    ANTENNAPARTIALMETALAREA 0.4356 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.924 LAYER METAL3 ;
    ANTENNAPARTIALMETALAREA 0.4356 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.924 LAYER METAL4 ;
  END i_in_data[20]
  PIN i_in_data[19] 
    ANTENNAPARTIALMETALAREA 81.7936 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 285.817 LAYER METAL2 ;
    ANTENNAPARTIALMETALAREA 0.4356 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.924 LAYER METAL3 ;
    ANTENNAPARTIALMETALAREA 0.4356 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.924 LAYER METAL4 ;
  END i_in_data[19]
  PIN i_in_data[18] 
    ANTENNAPARTIALMETALAREA 81.7186 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 285.415 LAYER METAL2 ;
    ANTENNAPARTIALMETALAREA 0.4356 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.924 LAYER METAL3 ;
    ANTENNAPARTIALMETALAREA 0.4356 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.924 LAYER METAL4 ;
  END i_in_data[18]
  PIN i_in_data[17] 
    ANTENNAPARTIALMETALAREA 15.4036 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 53.312 LAYER METAL3 ;
    ANTENNAPARTIALMETALAREA 0.4356 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.924 LAYER METAL4 ;
  END i_in_data[17]
  PIN i_in_data[16] 
    ANTENNAPARTIALMETALAREA 1.7676 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.586 LAYER METAL3 ;
    ANTENNAPARTIALMETALAREA 0.4356 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.924 LAYER METAL4 ;
  END i_in_data[16]
  PIN i_in_data[15] 
    ANTENNAPARTIALMETALAREA 14.692 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 51.422 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 71.49 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 250.355 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 37.008 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 129.808 LAYER METAL5 ;
  END i_in_data[15]
  PIN i_in_data[14] 
    ANTENNAPARTIALMETALAREA 15.06 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 52.71 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 64.848 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 227.108 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 35.352 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 124.012 LAYER METAL5 ;
  END i_in_data[14]
  PIN i_in_data[13] 
    ANTENNAPARTIALMETALAREA 0.198 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.693 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.96 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 51.326 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 180.061 LAYER METAL5 ;
  END i_in_data[13]
  PIN i_in_data[12] 
    ANTENNAPARTIALMETALAREA 15.796 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 55.286 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 45.25 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 158.515 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 35.168 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 123.368 LAYER METAL5 ;
  END i_in_data[12]
  PIN i_in_data[11] 
    ANTENNAPARTIALMETALAREA 50.012 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 175.042 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 32.066 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 112.371 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 1.162 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 4.207 LAYER METAL5 ;
  END i_in_data[11]
  PIN i_in_data[10] 
    ANTENNAPARTIALMETALAREA 50.206 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 175.721 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 20.2036 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 70.252 LAYER METAL4 ;
  END i_in_data[10]
  PIN i_in_data[9] 
    ANTENNAPARTIALMETALAREA 49.468 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 173.138 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 8.4576 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 29.141 LAYER METAL4 ;
  END i_in_data[9]
  PIN i_in_data[8] 
    ANTENNAPARTIALMETALAREA 19.292 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 67.522 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.304 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.204 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 29.958 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 104.993 LAYER METAL5 ;
  END i_in_data[8]
  PIN i_in_data[7] 
    ANTENNAPARTIALMETALAREA 21.132 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 73.962 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 10.81 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 37.975 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 75.612 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 264.782 LAYER METAL5 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA56 ;
    ANTENNAPARTIALMETALAREA 0.854 LAYER METAL6 ;
    ANTENNAPARTIALMETALSIDEAREA 3.269 LAYER METAL6 ;
  END i_in_data[7]
  PIN i_in_data[6] 
    ANTENNAPARTIALMETALAREA 20.948 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 73.318 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 19.748 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 69.258 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 84.302 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 295.197 LAYER METAL5 ;
  END i_in_data[6]
  PIN i_in_data[5] 
    ANTENNAPARTIALMETALAREA 76.24 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 266.84 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 28.44 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 99.68 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 24.53 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 85.995 LAYER METAL5 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA56 ;
    ANTENNAPARTIALMETALAREA 0.96 LAYER METAL6 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5 LAYER METAL6 ;
  END i_in_data[5]
  PIN i_in_data[4] 
    ANTENNAPARTIALMETALAREA 19.718 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 69.153 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.796 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.926 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 77.738 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 272.223 LAYER METAL5 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA56 ;
    ANTENNAPARTIALMETALAREA 0.632 LAYER METAL6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.352 LAYER METAL6 ;
  END i_in_data[4]
  PIN i_in_data[3] 
    ANTENNAPARTIALMETALAREA 50.1916 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 175.07 LAYER METAL3 ;
    ANTENNAPARTIALMETALAREA 0.4356 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.924 LAYER METAL4 ;
  END i_in_data[3]
  PIN i_in_data[2] 
    ANTENNAPARTIALMETALAREA 76.442 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 267.547 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 85.5936 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 299.117 LAYER METAL3 ;
    ANTENNAPARTIALMETALAREA 0.4356 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.924 LAYER METAL4 ;
  END i_in_data[2]
  PIN i_in_data[1] 
    ANTENNAPARTIALMETALAREA 0.5 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.75 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 73.8556 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 258.174 LAYER METAL3 ;
    ANTENNAPARTIALMETALAREA 0.4356 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.924 LAYER METAL4 ;
  END i_in_data[1]
  PIN i_in_data[0] 
    ANTENNAPARTIALMETALAREA 75.212 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 263.242 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 63.2496 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 220.913 LAYER METAL3 ;
    ANTENNAPARTIALMETALAREA 0.4356 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.924 LAYER METAL4 ;
  END i_in_data[0]
  PIN o_in_ready 
    ANTENNADIFFAREA 0.2176 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 16.357 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 57.3895 LAYER METAL2 ;
  END o_in_ready
  PIN o_out_valid 
    ANTENNADIFFAREA 0.413 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 16.347 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 57.3545 LAYER METAL2 ;
  END o_out_valid
  PIN o_out_data[23] 
    ANTENNAPARTIALMETALAREA 14.932 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 52.262 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 30.694 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 107.569 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.7208 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 42.124 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 147.574 LAYER METAL4 ;
  END o_out_data[23]
  PIN o_out_data[22] 
    ANTENNAPARTIALMETALAREA 15.424 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 53.984 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 20.206 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 70.861 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.7208 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 41.058 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 143.843 LAYER METAL4 ;
  END o_out_data[22]
  PIN o_out_data[21] 
    ANTENNAPARTIALMETALAREA 15.844 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 55.454 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 9.074 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 31.899 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.7208 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 45.588 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 159.698 LAYER METAL4 ;
  END o_out_data[21]
  PIN o_out_data[20] 
    ANTENNAPARTIALMETALAREA 15.178 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 53.123 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 2.266 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.071 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.7208 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 41.386 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 144.991 LAYER METAL4 ;
  END o_out_data[20]
  PIN o_out_data[19] 
    ANTENNAPARTIALMETALAREA 17.802 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 62.307 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 0.15 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER METAL5 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA56 ;
    ANTENNADIFFAREA 0.7208 LAYER METAL6 ; 
    ANTENNAPARTIALMETALAREA 37.778 LAYER METAL6 ;
    ANTENNAPARTIALMETALSIDEAREA 132.363 LAYER METAL6 ;
  END o_out_data[19]
  PIN o_out_data[18] 
    ANTENNAPARTIALMETALAREA 18.048 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 63.168 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.518 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.953 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 0.334 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.309 LAYER METAL5 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA56 ;
    ANTENNADIFFAREA 0.7208 LAYER METAL6 ; 
    ANTENNAPARTIALMETALAREA 31.874 LAYER METAL6 ;
    ANTENNAPARTIALMETALSIDEAREA 111.699 LAYER METAL6 ;
  END o_out_data[18]
  PIN o_out_data[17] 
    ANTENNAPARTIALMETALAREA 19.278 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 67.473 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.144 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 0.242 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.987 LAYER METAL5 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA56 ;
    ANTENNADIFFAREA 0.7208 LAYER METAL6 ; 
    ANTENNAPARTIALMETALAREA 30.152 LAYER METAL6 ;
    ANTENNAPARTIALMETALSIDEAREA 105.672 LAYER METAL6 ;
  END o_out_data[17]
  PIN o_out_data[16] 
    ANTENNADIFFAREA 0.7208 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 55.252 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 193.522 LAYER METAL2 ;
  END o_out_data[16]
  PIN o_out_data[15] 
    ANTENNADIFFAREA 0.5776 LAYER METAL2 ; 
    ANTENNAPARTIALMETALAREA 60.116 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 210.686 LAYER METAL2 ;
  END o_out_data[15]
  PIN o_out_data[14] 
    ANTENNAPARTIALMETALAREA 51.227 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 179.294 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 48.634 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 170.359 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.5776 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 11.138 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 39.123 LAYER METAL4 ;
  END o_out_data[14]
  PIN o_out_data[13] 
    ANTENNAPARTIALMETALAREA 55.908 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 195.678 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.5776 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 63.034 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 220.759 LAYER METAL4 ;
  END o_out_data[13]
  PIN o_out_data[12] 
    ANTENNAPARTIALMETALAREA 2.823 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.8805 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.5776 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 36.452 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 127.862 LAYER METAL4 ;
  END o_out_data[12]
  PIN o_out_data[11] 
    ANTENNAPARTIALMETALAREA 56.644 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 198.254 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.5776 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 45.3 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 158.69 LAYER METAL4 ;
  END o_out_data[11]
  PIN o_out_data[10] 
    ANTENNAPARTIALMETALAREA 51.724 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 181.174 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.7208 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 12.204 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 42.854 LAYER METAL4 ;
  END o_out_data[10]
  PIN o_out_data[9] 
    ANTENNAPARTIALMETALAREA 55.302 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 193.697 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.7208 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 12.88 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 45.22 LAYER METAL4 ;
  END o_out_data[9]
  PIN o_out_data[8] 
    ANTENNAPARTIALMETALAREA 56.256 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 196.896 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.7208 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 14.5 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 50.89 LAYER METAL4 ;
  END o_out_data[8]
  PIN o_out_data[7] 
    ANTENNADIFFAREA 0.7208 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 40.694 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 142.569 LAYER METAL3 ;
  END o_out_data[7]
  PIN o_out_data[6] 
    ANTENNADIFFAREA 0.7208 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 40.03 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 140.105 LAYER METAL3 ;
  END o_out_data[6]
  PIN o_out_data[5] 
    ANTENNAPARTIALMETALAREA 41.798 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 146.433 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.7208 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 4.814 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 16.989 LAYER METAL4 ;
  END o_out_data[5]
  PIN o_out_data[4] 
    ANTENNADIFFAREA 0.7208 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 40.132 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 140.602 LAYER METAL3 ;
  END o_out_data[4]
  PIN o_out_data[3] 
    ANTENNADIFFAREA 0.7208 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 36.912 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 129.332 LAYER METAL3 ;
  END o_out_data[3]
  PIN o_out_data[2] 
    ANTENNADIFFAREA 0.7208 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 37.372 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 130.942 LAYER METAL3 ;
  END o_out_data[2]
  PIN o_out_data[1] 
    ANTENNAPARTIALMETALAREA 2.732 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.562 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.7208 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 20.814 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 72.989 LAYER METAL4 ;
  END o_out_data[1]
  PIN o_out_data[0] 
    ANTENNADIFFAREA 0.7208 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 36.452 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 127.722 LAYER METAL3 ;
  END o_out_data[0]
END ipdc

END LIBRARY
