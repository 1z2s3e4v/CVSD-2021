/home/raid7_1/userd/d10013/CVSD/hw5/sram_lef/sram_256x8_ant.lef