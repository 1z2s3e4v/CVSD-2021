/home/raid7_1/userd/d10013/CVSD/lab6/Lab6/library/lef/antenna_8.lef