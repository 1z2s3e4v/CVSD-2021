/home/raid7_1/userd/d10013/CVSD/hw5/APR/library/lef/antenna_8.lef