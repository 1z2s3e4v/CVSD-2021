/home/raid7_1/userd/d10013/CVSD/hw5/APR/library/lef/tsmc13fsg_8lm_cic.lef